module foo();

initial
begin
  $display("hello world !!");
end

endmodule
